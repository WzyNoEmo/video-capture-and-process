
`timescale 1 ns / 1 ps

module GTP_DRM18K_WRAPPER
#(
    parameter [2:0] CSA_MASK = 3'b000,
    parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 18, // 1 2 4 8 16 32 9 18 36
    parameter integer DATA_WIDTH_B = 18, // 1 2 4 8 16 32 9 18 36
    parameter WRITE_MODE_A = "NORMAL_WRITE", // TRANSPARENT_WRITE READ_BEFORE_WRITE
    parameter WRITE_MODE_B = "NORMAL_WRITE", // TRANSPARENT_WRITE READ_BEFORE_WRITE
    parameter OUTPUT_REG_A = 0,
    parameter OUTPUT_REG_B = 0,
    parameter RESET_TYPE = "SYNC_RESET", // ASYNC_RESET ASYNC_RESET_SYNC_RELEASE

    parameter RAM_MODE = "TRUE_DUAL_PORT",  // SIMPLE_DUAL_PORT SINGLE_PORT ROM
    parameter WRITE_COLLISION_ARBITER = "NULL", // PORTA PORTB
    parameter GRS_EN = "TRUE",             //"TRUE"; "FALSE"
    parameter CLKA_OR_POL_INV = 1'b0,   //clka polarity invert for output register
    parameter CLKB_OR_POL_INV = 1'b0,   //clkb polarity invert for output register
    parameter INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
//add for initialization memory
    parameter BLOCK_X = 0         , //indicate X location of block memory when cascaded with DRM18Ks
    parameter BLOCK_Y = 0         , //indicate Y location of block memory when cascaded with DRM18Ks
    parameter RAM_DATA_WIDTH = 9  , //the total DATA WIDTH of cascaded DRMS
    parameter RAM_ADDR_WIDTH = 11 , //the total ADDR WIDTH of cascaded DRMS
    parameter INIT_FORMAT = "BIN"   //initial file data type binary or hexadecimal
) (
    output [17:0] QA,
    input [13:0] ADA,
    input ADAS,
    input [17:0] DA,
    input [2:0] CSA,
    input WEA,
    input CLKA, CEA, OCEA, RSTA,

    output [17:0] QB,
    input [13:0] ADB,
    input ADBS,
    input [17:0] DB,
    input [2:0] CSB,
    input WEB,
    input CLKB, CEB, OCEB, RSTB,
    output WWCONF
);

    GTP_DRM18K #(
    .GRS_EN(GRS_EN),
    .CSA_MASK(CSA_MASK),
    .CSB_MASK(CSB_MASK),
    .DATA_WIDTH_A(DATA_WIDTH_A),
    .DATA_WIDTH_B(DATA_WIDTH_B),
    .WRITE_MODE_A(WRITE_MODE_A),
    .WRITE_MODE_B(WRITE_MODE_B),
    .DOA_REG(OUTPUT_REG_A),
    .DOB_REG(OUTPUT_REG_B),
    .DOA_REG_CLKINV(CLKA_OR_POL_INV),
    .DOB_REG_CLKINV(CLKB_OR_POL_INV),
    .RST_TYPE( (RESET_TYPE == "SYNC_RESET") ? "SYNC" : ((RESET_TYPE == "ASYNC_RESET") ?  "ASYNC" : "ASYNC_SYNC_RELEASE") ),
    .RAM_MODE(RAM_MODE),
    .WRITE_COLLISION_ARBITER(WRITE_COLLISION_ARBITER),
    .INIT_00(INIT_00),
    .INIT_01(INIT_01),
    .INIT_02(INIT_02),
    .INIT_03(INIT_03),
    .INIT_04(INIT_04),
    .INIT_05(INIT_05),
    .INIT_06(INIT_06),
    .INIT_07(INIT_07),
    .INIT_08(INIT_08),
    .INIT_09(INIT_09),
    .INIT_0A(INIT_0A),
    .INIT_0B(INIT_0B),
    .INIT_0C(INIT_0C),
    .INIT_0D(INIT_0D),
    .INIT_0E(INIT_0E),
    .INIT_0F(INIT_0F),
    .INIT_10(INIT_10),
    .INIT_11(INIT_11),
    .INIT_12(INIT_12),
    .INIT_13(INIT_13),
    .INIT_14(INIT_14),
    .INIT_15(INIT_15),
    .INIT_16(INIT_16),
    .INIT_17(INIT_17),
    .INIT_18(INIT_18),
    .INIT_19(INIT_19),
    .INIT_1A(INIT_1A),
    .INIT_1B(INIT_1B),
    .INIT_1C(INIT_1C),
    .INIT_1D(INIT_1D),
    .INIT_1E(INIT_1E),
    .INIT_1F(INIT_1F),
    .INIT_20(INIT_20),
    .INIT_21(INIT_21),
    .INIT_22(INIT_22),
    .INIT_23(INIT_23),
    .INIT_24(INIT_24),
    .INIT_25(INIT_25),
    .INIT_26(INIT_26),
    .INIT_27(INIT_27),
    .INIT_28(INIT_28),
    .INIT_29(INIT_29),
    .INIT_2A(INIT_2A),
    .INIT_2B(INIT_2B),
    .INIT_2C(INIT_2C),
    .INIT_2D(INIT_2D),
    .INIT_2E(INIT_2E),
    .INIT_2F(INIT_2F),
    .INIT_30(INIT_30),
    .INIT_31(INIT_31),
    .INIT_32(INIT_32),
    .INIT_33(INIT_33),
    .INIT_34(INIT_34),
    .INIT_35(INIT_35),
    .INIT_36(INIT_36),
    .INIT_37(INIT_37),
    .INIT_38(INIT_38),
    .INIT_39(INIT_39),
    .INIT_3A(INIT_3A),
    .INIT_3B(INIT_3B),
    .INIT_3C(INIT_3C),
    .INIT_3D(INIT_3D),
    .INIT_3E(INIT_3E),
    .INIT_3F(INIT_3F),
    .INIT_FILE(INIT_FILE),
    .BLOCK_X(BLOCK_X),
    .BLOCK_Y(BLOCK_Y),
    .RAM_DATA_WIDTH(RAM_DATA_WIDTH),
    .RAM_ADDR_WIDTH(RAM_ADDR_WIDTH),
    .INIT_FORMAT(INIT_FORMAT)
    ) drm18k (
    .DOA(QA),
    .DOB(QB),
    .WWCONF(WWCONF),
    .DIA(DA),
    .DIB(DB),
    .ADDRA(ADA),
    .ADDRA_HOLD(ADAS),
    .ADDRB(ADB),
    .ADDRB_HOLD(ADBS),
    .CSA(CSA),
    .CSB(CSB),
    .CLKA(CLKA),
    .CLKB(CLKB),
    .CEA(CEA),
    .CEB(CEB),
    .WEA(WEA),
    .WEB(WEB),
    .ORCEA(OCEA),
    .ORCEB(OCEB),
    .RSTA(RSTA),
    .RSTB(RSTB)
    );

endmodule
